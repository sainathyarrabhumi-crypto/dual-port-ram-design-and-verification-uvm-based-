package ram_test_pkg;


//import uvm_pkg.sv
	import uvm_pkg::*;
//include uvm_macros.sv
	`include "uvm_macros.svh"
`include "tb_defs.sv"
`include "write_xtn.sv"
`include "ram_wr_agent_config.sv"
`include "ram_rd_agent_config.sv"
`include "ram_env_config.sv"
`include "ram_wr_driver.sv"
`include "ram_wr_monitor.sv"
`include "ram_wr_sequencer.sv"
`include "ram_wr_agent.sv"
`include "ram_wr_agt_top.sv"
`include "ram_wr_seqs.sv"

`include "read_xtn.sv"
`include "ram_rd_monitor.sv"
`include "ram_rd_sequencer.sv"
`include "ram_rd_seqs.sv"
`include "ram_rd_driver.sv"
`include "ram_rd_agent.sv"
`include "ram_rd_agt_top.sv"

`include "ram_virtual_sequencer.sv"
`include "ram_virtual_seqs.sv"
`include "ram_scoreboard.sv"

`include "ram_tb.sv"


`include "ram_vtest_lib.sv"
endpackage
